library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
USE ieee.numeric_std.all;


entity FSM_control24 is
  port( clock_25Mhz, v_sync, done, run	: in std_logic;
		x_t 		: out std_logic_vector(9 downto 1);
		y_t			: out std_logic_vector(8 downto 1);
		start		: out std_logic;
		color		: out std_logic_vector(2 downto 0));
		
end FSM_control24;

architecture seq of FSM_control24 is
  -- State definition:
  type states is (s0,ss0,s1, s2, s3, s4, s5, swb, swsquare, swait);
  
  signal st : states := s0;
  signal x_new : std_logic_vector(9 downto 1) := "000000000";
  signal x_old : std_logic_vector(9 downto 1) := "000000000";
  signal y_new : std_logic_vector(8 downto 1) := "00000000";
  signal y_old : std_logic_vector(8 downto 1) := "00000000";
  
  signal ld_col, ld_x, CE_new, sel_x, sel_col, ld_old : std_logic := '0';
  
  

begin

	--y_t <= "01000000";  -- VALUE = 64
	process(clock_25Mhz)
	Begin
		if (clock_25Mhz'event and clock_25Mhz='1') then
			case st is
				when s0 =>
					if(run = '1') then 
						st <= ss0;
					end if;
				when ss0 =>
					if(v_sync='0') then
						st <= s1;
					end if;
				when s1	=>
					st <= s2;
				when s2 =>
					st <= swb;
				when swb =>
					if(done='1') then		-- already erased
						st <= s3;
					end if;
				when s3 =>
					st <= s4;
				when s4 =>
					st <= s5;
				when s5 =>
					st <= swsquare;
				when swsquare =>	
					if(done='1') then		-- already drawn
						st <= swait;
					end if;
				when swait =>
					if(v_sync='1') then
						st <= s0;
					end if;
			End Case;
		End If;
	End Process;
	
		
	
-- Control signals generated by the control unit
--------
ld_x <= '1' when st=s1 or st=s4 else '0';
ld_col <= '1' when st=s1 or st=s4 else '0';
CE_new <= '1' when st=s1 else '0';
start <= '1' when st=s2 or st=s5 else '0';
ld_old <= '1' when st=s4 else '0';
sel_x <= '1' when st=s3 else '0' when st=ss0;
sel_col <= '1' when st=s3 else '0' when st=ss0;

	process(clock_25Mhz)
		Begin
			if (clock_25Mhz'event and clock_25Mhz='1') then
				-- color_t is the output of a register. Only two possible output values
				if ld_col = '1' and sel_col = '1' then
					color <= "010";
				elsif ld_col = '1' then
					color <= "000";
				end if;
				
				-- x_old
				if ld_old= '1' then
					x_old <= x_new;
					y_old <= y_new;
				end if;
				
				-- x_new
				if CE_new = '1' and x_new < "101000000" then
					x_new <= x_new+2;
				elsif CE_new = '1' then
					x_new <="000000000";
				end if;
				-- y_new
				if CE_new = '1' and y_new < "11110000" then
					y_new <= y_new+2;
				elsif CE_new = '1' then
					y_new <="00000000";
				end if;
				
				if ld_x = '1' and sel_x = '1' then	
					x_t <= x_new;
					y_t <= y_new;
					
				elsif ld_x = '1' then
					x_t <= x_old;
					y_t <= y_old;
				end if;
				
			
			End If;
		End Process;


End;