---------------------------------------------------------------------------------------
-- code_v1: Main controller of design version 1:
-- Generates START signal when button(0) is pressed........................................................................................
-- Reades from switches and forms the bus x_t
-- Author: Pol Carrera and Marc Martinez. Date: 31-10-2019.
-- Electronic System Design for Communications - ESDC - ETSTB. UPC. Barcelona.
----------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;


entity code_v3 is
  port( clk_25          	: in std_logic;
		GO			        : out std_logic;
		sw, btn 		    : in std_logic_vector(3 downto 0) );
end code_v3;

architecture state_machine of code_v3 is
  -- State definition:
  type states is (wait_s0, s1, s2, wait_s3, s4, OK_s5, KO_s5, wait_s6, s7, OK_s8,
                  wait_s9, s10, s11, wait_s12, s13, OK_s14, KO_s14, wait_s15, s16, OK_s17);
  
  -- output of register state:
  signal st : states := wait_s0;

  Begin
 
 -- Control State Machine
 -- Description
    -- st<=wait_s0;
	process(clk_25)
	Begin
		if (clk_25'event and clk_25='1') then
			case st is
				when wait_s0 =>
					if(btn(0) = '1') then 
						st <= s1;
					end if;
				when s1 =>
					if(sw = "0001") then 
						st <= s2;
					else
					    st <= wait_s0;
				    end if;
				when s2 =>
					if(btn(0) = '0') then 
						st <= wait_s3;
					end if;
				when wait_s3 =>
					if(btn(0) = '1') then 
						st <= s4;
					end if;
				when s4 =>
					if(sw = "0011") then 
						st <= OK_s5;
					elsif(sw = "0001") then 
						st <= s2;
					else
					    st <= KO_s5;
				    end if;
				when KO_s5 =>
					if(btn(0) = '0') then 
						st <= wait_s0;
					end if;
			    when OK_s5 =>
					if(btn(0) = '0') then 
						st <= wait_s6;
					end if;
				when wait_s6 =>
					if(btn(0) = '1') then 
						st <= s7;
					end if;
				when s7 =>
					if(sw = "0111") then 
						st <= OK_s8;
					elsif(sw = "0001") then 
						st <= s2;
					else
					    st <= KO_s5;
				    end if;
				when OK_s8 =>
					if(btn(0) = '0') then 
						st <= wait_s9;
					end if;





				when wait_s9 =>
					if(btn(0) = '1') then 
						st <= s10;
					end if;
				when s10 =>
					if(sw = "0001") then 
						st <= s11;
					else
					    st <= wait_s9;
				    end if;
				when s11 =>
					if(btn(0) = '0') then 
						st <= wait_s12;
					end if;
				when wait_s12 =>
					if(btn(0) = '1') then 
						st <= s13;
					end if;
				when s13 =>
					if(sw = "0011") then 
						st <= OK_s14;
					elsif(sw = "0001") then 
						st <= s11;
					else
					    st <= KO_s14;
				    end if;
				when KO_s14 =>
					if(btn(0) = '0') then 
						st <= wait_s9;
					end if;
			    when OK_s14 =>
					if(btn(0) = '0') then 
						st <= wait_s15;
					end if;
				when wait_s15 =>
					if(btn(0) = '1') then 
						st <= s16;
					end if;
				when s16 =>
					if(sw = "0111") then 
						st <= OK_s17;
					elsif(sw = "0001") then 
						st <= s11;
					else
					    st <= KO_s14;
				    end if;
				when OK_s17 =>
					if(btn(0) = '0') then 
						st <= wait_s0;
					end if;

			End Case;
		End If;
	End Process;
	
-- Control signals generated by the control unit
GO <= '1' when st = wait_s9 or st=s10 or st=s11 or st=wait_s12 or st=s13 or st=KO_s14 or st=OK_s14 or st=wait_s15 or st=s16 or st=OK_s17 else '0';
			
End state_machine;
						
			
				
				
				